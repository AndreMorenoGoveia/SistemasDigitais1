`timescale 1ms/100ns

module testbench;

    wire [3:0] h1;
    wire [3:0] h2;
    wire [3:0] h3;
    wire [3:0] h4;

    main inst0 ();


endmodule